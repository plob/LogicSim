module c17 (N1,N2,N3,N20);

input N1,N2,N3;

output N20;

xor AND (N20, N1, N2, N3);

endmodule
